//================================================
//  University  : UIT - www.uit.edu.vn
//  Course name : System-on-Chip Design
//  Lab name    : lab3
//  File name   : rom.v
//  Author      : Pham Thanh Hung
//  Date        : Oct 21, 2017
//  Version     : 1.0
//-------------------------------------------------
// Modification History
//
//================================================
module rom(
//input
addr,
//output
data
);

input [31:0] addr;
output [31:0] data;

reg [31:0] data;
`define ADD 6'b100000
`define SUB 6'b100010
`define OP_0 6'h0
`define LW 6'b100011
//
//reg [31:0] mem [0:1023];
//assign data = mem[addr];
//op-6bit|rd-5bit|rt-5bit|rs-5bit|shamt-5bit|function-6bit|
//ADD R3,R2,R1;
//SUB R4,R3,R7;
//LW  R8,4(R3);

always @(*) begin
    case(addr)
//        //32'h00000000: data = 32'b00000001001010101010000000100000;
//        32'h00000000: data = {`OP_0,3,2,1,0,`ADD};
//        //32'h00000004: data = 32'b00000001001010101010000000100000;
//        32'h00000004: data = {`OP_0,4,3,7,0,`SUB};
//        //32'h00000008: data = 32'b00000001001010101010000000100000;
//        32'h00000008: data = {`LW,3,8,4};
//        32'h0000000c: data = 32'b00000001001010101010000000100000;
//        32'h00000010: data = 32'b00000001001010101010000000100000;
//        32'h00000014: data = 32'b10101111101001000000000000000000;
//        32'h00000018: data = 32'b10001111101010000000000000000000;
//        32'h0000001c: data = 32'b00010000001000000000000000000011;
        32'h00000000: data = 32'b00111100000000100000000000000101;
        32'h00000004: data = 32'b00111100000000110000000000001101;
        32'h00000008: data = 32'b00100000000001000000000000010011;
        32'h0000000c: data = 32'b00100000000001010000000000001100;
        32'h00000010: data = 32'b00100000000011011111111010011100;
        32'h00000014: data = 32'b00000000010000110000100000100000;
        32'h00000018: data = 32'b00000000011000100011000000100010;
        32'h0000001c: data = 32'b10101100101000110000000000000000;
        32'h00000020: data = 32'b00000000010000110011100000100100;
        32'h00000024: data = 32'b00000000010000110100000000100101;
        32'h00000028: data = 32'b00000000010000110100100000101010;
        32'h0000002c: data = 32'b00000001101000110110000000101010;
        32'h00000030: data = 32'b10001100101010100000000000000000;
        32'h00000034: data = 32'b10101100101000010000000000000000;
        32'h00000038: data = 32'b00100000000001000000000001111001;
        32'h0000003c: data = 32'b00010001010000110000000000000001;
        32'h00000040: data = 32'b00100000000010110000000000001111;
//        32'h00000038: data = ;
//        32'h0000003c: data = ;
        //insert your instructions here
        default: data = 32'hFFFF_FFFF;
    endcase

end

endmodule
